package jtag_agent_pkg ;
   import uvm_pkg::*;
   import jtag_def_pkg::*;
`include "uvm_macros.svh"

`include "jtag_agent_cfg.svh"
`include "jtag_transaction.svh"
`include "jtag_sequence_lib.svh"
`include "jtag_sequencer.svh"
`include "jtag_monitor.svh"
`include "jtag_driver.svh"
`include "jtag_agent.svh"

endpackage // pack_all
   