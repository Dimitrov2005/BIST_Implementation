package env_pkg ;
   import uvm_pkg::*;
   import def_pkg::*;
   
   import stac_agent_pkg::*;
`include "uvm_macros.svh"

`include "Scoreboard.svh"
`include "env_config.svh"
`include "Environment.svh"
`include "test.svh"

endpackage // pack_all
   