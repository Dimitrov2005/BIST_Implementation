package env_pkg ;
	import uvm_pkg::*;
	import jtag_def_pkg::*;
	 // fuse def pkg ??? 
	import jtag_agent_pkg::*;
	import fuse_agent_pkg::*;
	
	`include "uvm_macros.svh"
	`include "Scoreboard.svh"
	`include "env_config.svh"
	`include "Environment.svh"
	`include "test.svh"

endpackage // pack_all
   