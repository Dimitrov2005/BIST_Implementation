package fuse_agent_pkg ;
   import uvm_pkg::*;
   import fuse_def_pkg::*;
`include "uvm_macros.svh"

`include "fuse_agent_cfg.svh"
`include "fuse_transaction.svh"
`include "fuse_sequence_lib.svh"
`include "fuse_sequencer.svh"
`include "fuse_monitor.svh"
`include "fuse_driver.svh"
`include "fuse_agent.svh"

endpackage // pack_all
   