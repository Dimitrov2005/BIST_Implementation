package stac_agent_pkg ;
   import uvm_pkg::*;
   import stac_def_pkg::*;
`include "uvm_macros.svh"

`include "stac_agent_cfg.svh"
`include "stac_transaction.svh"
`include "stac_sequence_lib.svh"
`include "stac_sequencer.svh"
`include "stac_monitor.svh"
`include "stac_driver.svh"
`include "stac_agent.svh"

endpackage // pack_all
   