package fuse_def_pkg;

parameter SIZE_TDR1=17;
parameter ADDR_TDR1= 8'h45;
parameter DEF_VAL_TDR1=17'ha;
parameter RO_TDR1=0;
parameter SIZE_TDR2=33;
parameter ADDR_TDR2=8'h77;
parameter DEF_VAL_TDR2=33'ha;
parameter RO_TDR2=1;
   
endpackage // def_pkg
   
   